module segmentos_letras(

 input [3:0] bin, //entradas binarias
 
 output reg [6:0] seg //salidas para el display de 7 segmentos
 
);
 
 //logica de decodificacion para el display de 7 segmentos
 
 always @(bin) 
  begin
    case (bin)
 
     4'b0000: seg= 7'b0001100; //P correcto
     4'b0001: seg= 7'b1000000; //O correcto
     4'b0010: seg= 7'b1000111; //L correcto
     4'b0011: seg= 7'b1000000; //O correcto
     4'b0100: seg= 7'b0111111; //- correcto
     4'b0101: seg= 7'b0010010; //S correcto
     4'b0110: seg= 7'b1000000; //O correcto
     4'b0111: seg= 7'b1000111; //L correcto
     4'b1000: seg= 7'b0001000; //A correcto
     4'b1001: seg= 7'b0111111; //- correcto
     4'b1010: seg= 7'b1000110; //C correcto
     4'b1011: seg= 7'b1000000; //O correcto
     4'b1100: seg= 7'b0010010; //S correcto
     4'b1101: seg= 7'b0001000; //A correcto
     4'b1110: seg= 7'b0010010; //S correcto
     4'b1111: seg= 7'b1111111; // correcto
 
     default: seg= 7'b1111111; //default correcto
 
    endcase

 
 end


endmodule

 